`include "const.v"

module IF_ID (
        input wire [`INST_ADDR_WIDTH - 1:0] inst_addr,
        input wire [`INST_WIDTH - 1:0] inst
    );

endmodule
